//Subject:     CO project 2 - PC
//--------------------------------------------------------------------------------
//Version:     1
//--------------------------------------------------------------------------------
//Writer:      Luke
//----------------------------------------------
//Date:        2010/8/16
//----------------------------------------------
//Description: 
//--------------------------------------------------------------------------------

module PC(
    clk_i,
	rst_i,
	pc_in_i,
	pc_out_o,
	pc_write
	);
     
//I/O ports
input			pc_write;
input           clk_i;
input	        rst_i;
input  [32-1:0] pc_in_i;
output [32-1:0] pc_out_o;
 
//Internal Signals
reg    [32-1:0] pc_out_o;
 
//Parameter

    
//Main function
always @(posedge clk_i) begin
    if(~rst_i)
	    pc_out_o <= 0;
	else if(pc_write)
		pc_out_o <=pc_out_o;
	else
	    pc_out_o <= pc_in_i;
end

endmodule



                    
                    